
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity calculator is
    Port ( n1 : in  STD_LOGIC_VECTOR(3 downto 0);
           n2 : in  STD_LOGIC_VECTOR(3 downto 0);
			  ope : in  STD_LOGIC_VECTOR(3 downto 0);
           result : out  STD_LOGIC);
end calculator;

architecture Behavioral of calculator is
	
begin

end Behavioral;

